3e 2b 2b 2b 2b 2b 2b 2b 2b 5b 3c 2b 2b 2b 2b 2b 2b 2b 2b 2b 3e 2d 5d 3c 2e 00